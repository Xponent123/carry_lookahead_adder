.include TSMC_180nm.txt

.param SUPPLY=1.8
.global gnd vdd  

Vdd	vdd	gnd	'SUPPLY'

VA0 a0 gnd pulse 1.8  0 0 100p 100p 10n 20n
VA1 a1 gnd pulse 1.8 0  0 100p 100p 10n 20n
VA2 a2 gnd pulse 1.8 0  0 100p 100p 10n 40n
VA3 a3 gnd pulse 1.8  0 0 100p 100p 10n 40n

VB0 b0 gnd pulse 1.8 0  0 100p 100p 10n 80n
VB1 b1 gnd pulse 1.8  0 0 100p 100p 10n 40n
VB2 b2 gnd pulse 1.8  0 0 100p 100p 10n 20n
VB3 b3 gnd pulse 1.8 0  0 100p 100p 10n 20n

VC0 c0 gnd pulse 1.8 0  0 100p 100p 10n 40n


.option scale=0.09u

M1000 a_685_911# c0 vdd w_670_905# CMOSP w=8 l=2
+  ad=216 pd=102 as=4256 ps=2424
M1001 a_253_1351# a1 gnd Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=1784 ps=1484
M1002 gnd a_339_785# a_334_788# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1003 a_33_1351# a0 gnd Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=0 ps=0
M1004 a_381_1315# a1 gnd Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1005 a_685_1089# a_536_696# gnd Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=0 ps=0
M1006 a_821_1315# a3 gnd Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1007 a_593_639# a_542_639# s3 Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=32 ps=24
M1008 a_122_639# c0 vdd w_109_651# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1009 vdd a_116_696# a_346_1058# w_331_1052# CMOSP w=8 l=2
+  ad=0 pd=0 as=136 ps=66
M1010 vdd a_256_696# a_495_988# w_480_982# CMOSP w=8 l=2
+  ad=0 pd=0 as=160 ps=72
M1011 a_685_988# a_256_696# vdd w_670_982# CMOSP w=8 l=2
+  ad=160 pd=72 as=0 ps=0
M1012 a_698_827# a_696_771# a_678_771# w_667_821# CMOSP w=8 l=2
+  ad=80 pd=36 as=56 ps=30
M1013 a_350_1315# a1 gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1014 a_570_1315# a2 vdd w_557_1327# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1015 a_229_792# a_63_1351# gnd Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=0 ps=0
M1016 a_503_1351# a_473_1383# vdd w_458_1377# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1017 a_433_639# a_334_788# gnd Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1018 vdd a_63_1351# a_346_1121# w_331_1115# CMOSP w=8 l=2
+  ad=0 pd=0 as=80 ps=36
M1019 s0 c0 a_153_707# w_139_701# CMOSP w=8 l=2
+  ad=64 pd=32 as=64 ps=32
M1020 vdd a_396_696# a_685_1058# w_670_1052# CMOSP w=8 l=2
+  ad=0 pd=0 as=136 ps=66
M1021 a_313_707# a_256_696# s1 w_279_701# CMOSP w=8 l=2
+  ad=64 pd=32 as=64 ps=32
M1022 a_262_689# a_256_696# vdd w_249_701# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1023 a_339_785# a_369_785# gnd Gnd CMOSN w=4 l=2
+  ad=68 pd=50 as=0 ps=0
M1024 vdd a_130_1315# a_181_1383# w_147_1377# CMOSP w=8 l=2
+  ad=0 pd=0 as=64 ps=32
M1025 vdd a_570_1315# a_621_1383# w_587_1377# CMOSP w=8 l=2
+  ad=0 pd=0 as=64 ps=32
M1026 a_495_988# a_396_696# vdd w_480_982# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1027 vdd a_396_696# a_685_988# w_670_982# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1028 a_495_1019# a_396_696# gnd Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=0 ps=0
M1029 vdd a_678_771# c4 w_667_821# CMOSP w=8 l=2
+  ad=0 pd=0 as=40 ps=26
M1030 a_253_1383# a1 vdd w_238_1377# CMOSP w=8 l=2
+  ad=80 pd=36 as=0 ps=0
M1031 vdd a_503_1351# a_685_1121# w_670_1115# CMOSP w=8 l=2
+  ad=0 pd=0 as=80 ps=36
M1032 a_346_1121# a_63_1351# a_346_1089# Gnd CMOSN w=4 l=2
+  ad=28 pd=22 as=40 ps=28
M1033 a_346_1019# a_256_696# gnd Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=0 ps=0
M1034 a_732_771# a_685_988# vdd w_670_982# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1035 a_253_1383# b1 a_253_1351# Gnd CMOSN w=4 l=2
+  ad=28 pd=22 as=0 ps=0
M1036 a_693_1383# b3 a_693_1351# Gnd CMOSN w=4 l=2
+  ad=28 pd=22 as=40 ps=28
M1037 gnd a_542_778# a_488_778# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=80 ps=56
M1038 gnd a_229_792# a_224_795# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1039 a_381_1383# a_350_1365# vdd w_367_1377# CMOSP w=8 l=2
+  ad=64 pd=32 as=0 ps=0
M1040 a_33_1383# a0 vdd w_18_1377# CMOSP w=8 l=2
+  ad=80 pd=36 as=0 ps=0
M1041 a_821_1383# a_790_1365# vdd w_807_1377# CMOSP w=8 l=2
+  ad=64 pd=32 as=0 ps=0
M1042 gnd a_720_771# a_678_771# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=108 ps=78
M1043 a_520_827# a_518_778# a_508_827# w_477_821# CMOSP w=8 l=2
+  ad=80 pd=36 as=80 ps=36
M1044 gnd a_402_689# a_453_639# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1045 a_130_1365# b0 gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1046 a_33_1383# b0 a_33_1351# Gnd CMOSN w=4 l=2
+  ad=28 pd=22 as=0 ps=0
M1047 a_790_1365# b3 gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1048 a_350_1365# b1 vdd w_337_1377# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1049 a_685_1121# a_503_1351# a_685_1089# Gnd CMOSN w=4 l=2
+  ad=28 pd=22 as=0 ps=0
M1050 a_685_1019# a_536_696# gnd Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=0 ps=0
M1051 a_369_785# a_346_1121# vdd w_331_1115# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1052 a_685_858# a_536_696# gnd Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=0 ps=0
M1053 a_346_1058# c0 vdd w_331_1052# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1054 a_153_639# c0 gnd Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1055 a_181_1315# a_130_1315# a_116_696# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=32 ps=24
M1056 a_621_1315# a_570_1315# a_396_696# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=32 ps=24
M1057 s1 a_256_696# a_293_639# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=32 ps=24
M1058 a_593_707# a_536_696# s3 w_559_701# CMOSP w=8 l=2
+  ad=64 pd=32 as=64 ps=32
M1059 a_685_911# a_536_696# vdd w_670_905# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1060 a_495_988# a_116_696# vdd w_480_982# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1061 vdd a_63_1351# a_685_988# w_670_982# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1062 a_402_639# a_334_788# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1063 a_369_785# a_346_1121# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1064 a_542_689# a_536_696# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1065 a_433_707# a_402_689# vdd w_419_701# CMOSP w=8 l=2
+  ad=64 pd=32 as=0 ps=0
M1066 gnd a_259_792# a_229_792# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1067 a_249_827# a_63_1351# a_229_792# w_218_821# CMOSP w=8 l=2
+  ad=80 pd=36 as=56 ps=30
M1068 a_283_1351# a_253_1383# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1069 a_236_1121# a_116_696# vdd w_221_1115# CMOSP w=8 l=2
+  ad=80 pd=36 as=0 ps=0
M1070 a_696_771# a_693_1383# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1071 vdd b1 a_253_1383# w_238_1377# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1072 vdd b3 a_693_1383# w_678_1377# CMOSP w=8 l=2
+  ad=0 pd=0 as=80 ps=36
M1073 a_358_1019# a_116_696# a_346_1019# Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=0 ps=0
M1074 a_63_1351# a_33_1383# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1075 gnd a_790_1365# a_841_1315# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1076 a_236_1089# a_116_696# gnd Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=0 ps=0
M1077 gnd a_122_689# a_173_639# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1078 a_381_785# a_346_1058# vdd w_331_1052# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1079 a_685_942# a_536_696# gnd Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=0 ps=0
M1080 vdd a_488_778# a_483_781# w_477_821# CMOSP w=8 l=2
+  ad=0 pd=0 as=40 ps=26
M1081 vdd b0 a_33_1383# w_18_1377# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1082 a_473_1351# a2 gnd Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=0 ps=0
M1083 a_488_778# a_503_1351# gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1084 a_709_858# a_256_696# a_697_858# Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=40 ps=28
M1085 a_542_778# a_495_988# vdd w_480_982# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1086 s3 a_536_696# a_573_639# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1087 vdd a_229_792# a_224_795# w_218_821# CMOSP w=8 l=2
+  ad=0 pd=0 as=40 ps=26
M1088 a_181_1383# b0 a_116_696# w_147_1377# CMOSP w=8 l=2
+  ad=0 pd=0 as=64 ps=32
M1089 a_621_1383# b2 a_396_696# w_587_1377# CMOSP w=8 l=2
+  ad=0 pd=0 as=64 ps=32
M1090 a_697_1019# a_396_696# a_685_1019# Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=0 ps=0
M1091 vdd a_381_785# a_371_827# w_328_821# CMOSP w=8 l=2
+  ad=0 pd=0 as=80 ps=36
M1092 a_122_639# c0 gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1093 a_678_771# a_732_771# gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1094 a_685_911# a_256_696# vdd w_670_905# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1095 a_601_1315# a2 gnd Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1096 vdd a_402_639# a_453_707# w_419_701# CMOSP w=8 l=2
+  ad=0 pd=0 as=64 ps=32
M1097 vdd a_256_696# a_495_1058# w_480_1052# CMOSP w=8 l=2
+  ad=0 pd=0 as=136 ps=66
M1098 a_262_689# a_256_696# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1099 a_153_707# a_122_689# vdd w_139_701# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1100 a_697_858# a_396_696# a_685_858# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1101 a_570_1315# a2 gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1102 s1 a_224_795# a_293_707# w_279_701# CMOSP w=8 l=2
+  ad=0 pd=0 as=64 ps=32
M1103 a_130_1315# a0 vdd w_117_1327# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1104 a_283_1351# a_253_1383# vdd w_238_1377# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1105 a_790_1315# a3 vdd w_777_1327# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1106 a_696_771# a_693_1383# vdd w_678_1377# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1107 a_402_689# a_396_696# vdd w_389_701# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1108 vdd a_396_696# a_685_911# w_670_905# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1109 vdd c0 a_236_1121# w_221_1115# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1110 vdd a_283_1351# a_495_1121# w_480_1115# CMOSP w=8 l=2
+  ad=0 pd=0 as=80 ps=36
M1111 vdd c0 a_495_988# w_480_982# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1112 a_722_827# a_720_771# a_710_827# w_667_821# CMOSP w=8 l=2
+  ad=80 pd=36 as=80 ps=36
M1113 a_63_1351# a_33_1383# vdd w_18_1377# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1114 vdd a_790_1315# a_841_1383# w_807_1377# CMOSP w=8 l=2
+  ad=0 pd=0 as=64 ps=32
M1115 a_507_942# a_256_696# a_495_942# Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=40 ps=28
M1116 a_709_942# a_256_696# a_697_942# Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=40 ps=28
M1117 vdd a_259_792# a_249_827# w_218_821# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1118 a_346_1058# c0 a_358_1019# Gnd CMOSN w=4 l=2
+  ad=28 pd=22 as=0 ps=0
M1119 a_116_696# b0 a_161_1315# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1120 a_396_696# b2 a_601_1315# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1121 a_473_1383# a2 vdd w_458_1377# CMOSP w=8 l=2
+  ad=80 pd=36 as=0 ps=0
M1122 a_236_1121# c0 a_236_1089# Gnd CMOSN w=4 l=2
+  ad=28 pd=22 as=0 ps=0
M1123 a_495_1121# a_283_1351# a_495_1089# Gnd CMOSN w=4 l=2
+  ad=28 pd=22 as=40 ps=28
M1124 a_542_639# a_483_781# vdd w_529_651# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1125 a_453_639# a_402_639# s2 Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1126 a_473_1383# b2 a_473_1351# Gnd CMOSN w=4 l=2
+  ad=28 pd=22 as=0 ps=0
M1127 gnd a_542_689# a_593_639# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1128 vdd a_122_639# a_173_707# w_139_701# CMOSP w=8 l=2
+  ad=0 pd=0 as=64 ps=32
M1129 a_601_1383# a_570_1365# vdd w_587_1377# CMOSP w=8 l=2
+  ad=64 pd=32 as=0 ps=0
M1130 a_495_942# a_396_696# gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1131 a_697_942# a_396_696# a_685_942# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1132 gnd a_518_778# a_488_778# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1133 a_721_858# a_116_696# a_709_858# Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=0 ps=0
M1134 a_350_1365# b1 gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1135 s3 a_483_781# a_573_707# w_559_701# CMOSP w=8 l=2
+  ad=0 pd=0 as=64 ps=32
M1136 a_570_1365# b2 vdd w_557_1377# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1137 a_259_792# a_236_1121# vdd w_221_1115# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1138 a_518_778# a_495_1121# vdd w_480_1115# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1139 a_495_1058# a_63_1351# vdd w_480_1052# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1140 a_401_1315# a_350_1315# a_256_696# Gnd CMOSN w=4 l=2
+  ad=32 pd=24 as=32 ps=24
M1141 a_732_771# a_685_988# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1142 a_122_689# a_116_696# vdd w_109_701# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1143 gnd a_744_771# a_678_771# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1144 vdd a_116_696# a_685_911# w_670_905# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1145 a_841_1315# a_790_1315# a_536_696# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1146 gnd a_381_785# a_339_785# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1147 a_381_785# a_346_1058# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1148 a_259_792# a_236_1121# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1149 a_518_778# a_495_1121# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1150 a_116_696# a0 a_161_1383# w_147_1377# CMOSP w=8 l=2
+  ad=0 pd=0 as=64 ps=32
M1151 a_396_696# a2 a_601_1383# w_587_1377# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1152 a_708_771# a_685_1121# vdd w_670_1115# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1153 a_685_1058# a_283_1351# vdd w_670_1052# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1154 a_262_639# a_224_795# vdd w_249_651# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1155 a_173_639# a_122_639# s0 Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1156 gnd a_262_689# a_313_639# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=32 ps=24
M1157 a_532_827# a_530_778# a_520_827# w_477_821# CMOSP w=8 l=2
+  ad=80 pd=36 as=0 ps=0
M1158 vdd b2 a_473_1383# w_458_1377# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1159 a_734_827# a_732_771# a_722_827# w_667_821# CMOSP w=8 l=2
+  ad=80 pd=36 as=0 ps=0
M1160 a_744_771# a_685_911# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1161 a_507_1019# a_256_696# a_495_1019# Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=0 ps=0
M1162 a_519_942# a_116_696# a_507_942# Gnd CMOSN w=4 l=2
+  ad=40 pd=28 as=0 ps=0
M1163 a_685_988# a_63_1351# a_709_942# Gnd CMOSN w=4 l=2
+  ad=28 pd=22 as=0 ps=0
M1164 a_708_771# a_685_1121# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1165 a_573_639# a_483_781# gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1166 gnd a_350_1365# a_401_1315# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1167 a_744_771# a_685_911# vdd w_670_905# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1168 a_530_778# a_495_1058# vdd w_480_1052# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1169 a_693_1351# a3 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1170 a_453_707# a_396_696# s2 w_419_701# CMOSP w=8 l=2
+  ad=0 pd=0 as=64 ps=32
M1171 gnd a_488_778# a_483_781# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1172 vdd a_542_639# a_593_707# w_559_701# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1173 a_401_1383# b1 a_256_696# w_367_1377# CMOSP w=8 l=2
+  ad=64 pd=32 as=64 ps=32
M1174 a_841_1383# b3 a_536_696# w_807_1377# CMOSP w=8 l=2
+  ad=0 pd=0 as=64 ps=32
M1175 a_402_689# a_396_696# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1176 a_161_1315# a0 gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1177 a_720_771# a_685_1058# vdd w_670_1052# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1178 a_678_771# a_708_771# gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1179 a_359_827# a_283_1351# a_339_785# w_328_821# CMOSP w=8 l=2
+  ad=80 pd=36 as=56 ps=30
M1180 a_790_1315# a3 gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1181 a_130_1315# a0 gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1182 a_542_778# a_495_988# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1183 a_350_1315# a1 vdd w_337_1327# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1184 a_293_639# a_224_795# gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1185 vdd a_350_1315# a_401_1383# w_367_1377# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1186 s2 a_396_696# a_433_639# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1187 gnd a_696_771# a_678_771# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1188 a_256_696# b1 a_381_1315# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1189 a_495_1058# a_63_1351# a_507_1019# Gnd CMOSN w=4 l=2
+  ad=28 pd=22 as=0 ps=0
M1190 a_542_639# a_483_781# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1191 a_536_696# b3 a_821_1315# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1192 a_173_707# a_116_696# s0 w_139_701# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1193 a_693_1383# a3 vdd w_678_1377# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1194 vdd a_262_639# a_313_707# w_279_701# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1195 vdd a_339_785# a_334_788# w_328_821# CMOSP w=8 l=2
+  ad=0 pd=0 as=40 ps=26
M1196 vdd a_744_771# a_734_827# w_667_821# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1197 vdd a_542_778# a_532_827# w_477_821# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1198 a_495_988# c0 a_519_942# Gnd CMOSN w=4 l=2
+  ad=28 pd=22 as=0 ps=0
M1199 a_573_707# a_542_689# vdd w_559_701# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1200 a_122_689# a_116_696# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1201 a_161_1383# a_130_1365# vdd w_147_1377# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1202 a_570_1365# b2 gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1203 a_685_1058# a_283_1351# a_697_1019# Gnd CMOSN w=4 l=2
+  ad=28 pd=22 as=0 ps=0
M1204 a_790_1365# b3 vdd w_777_1377# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1205 a_130_1365# b0 vdd w_117_1377# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1206 gnd a_678_771# c4 Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1207 a_495_1058# a_396_696# vdd w_480_1052# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1208 a_346_1058# a_256_696# vdd w_331_1052# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1209 a_530_778# a_495_1058# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1210 s0 a_116_696# a_153_639# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1211 a_402_639# a_334_788# vdd w_389_651# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1212 a_371_827# a_369_785# a_359_827# w_328_821# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1213 gnd a_283_1351# a_339_785# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1214 a_256_696# a1 a_381_1383# w_367_1377# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1215 a_495_1121# a_396_696# vdd w_480_1115# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1216 a_685_988# a_536_696# vdd w_670_982# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1217 a_313_639# a_262_639# s1 Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1218 a_262_639# a_224_795# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1219 a_536_696# a3 a_821_1383# w_807_1377# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1220 a_346_1121# a_256_696# vdd w_331_1115# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1221 a_503_1351# a_473_1383# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1222 a_685_1058# a_536_696# vdd w_670_1052# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1223 a_293_707# a_262_689# vdd w_279_701# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1224 a_720_771# a_685_1058# gnd Gnd CMOSN w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1225 s2 a_334_788# a_433_707# w_419_701# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1226 a_495_1089# a_396_696# gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1227 a_488_778# a_530_778# gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1228 a_685_911# c0 a_721_858# Gnd CMOSN w=4 l=2
+  ad=28 pd=22 as=0 ps=0
M1229 gnd a_130_1365# a_181_1315# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1230 gnd a_570_1365# a_621_1315# Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1231 a_346_1089# a_256_696# gnd Gnd CMOSN w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1232 a_542_689# a_536_696# vdd w_529_701# CMOSP w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1233 a_685_1121# a_536_696# vdd w_670_1115# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1234 a_710_827# a_708_771# a_698_827# w_667_821# CMOSP w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1235 a_508_827# a_503_1351# a_488_778# w_477_821# CMOSP w=8 l=2
+  ad=0 pd=0 as=56 ps=30
C0 a_369_785# a_381_785# 0.85fF
C1 a_116_696# a_63_1351# 7.59fF
C2 w_18_1377# a_63_1351# 0.03fF
C3 a_130_1315# gnd 0.31fF
C4 a_262_689# a_262_639# 0.02fF
C5 vdd w_117_1377# 0.05fF
C6 a_283_1351# w_328_821# 0.06fF
C7 a_122_689# vdd 0.74fF
C8 a_63_1351# a_259_792# 0.99fF
C9 a_381_785# w_328_821# 0.06fF
C10 w_419_701# a_402_639# 0.06fF
C11 a_685_988# a_732_771# 0.05fF
C12 a_350_1315# gnd 0.31fF
C13 w_807_1377# vdd 0.11fF
C14 vdd a_542_689# 0.74fF
C15 vdd w_557_1377# 0.05fF
C16 w_367_1377# a_256_696# 0.02fF
C17 w_670_982# a_536_696# 0.06fF
C18 w_367_1377# b1 0.06fF
C19 vdd a_685_911# 0.21fF
C20 a_130_1365# a_116_696# 0.08fF
C21 vdd w_559_701# 0.11fF
C22 w_218_821# a_63_1351# 0.06fF
C23 a_253_1383# gnd 0.04fF
C24 w_559_701# a_542_689# 0.19fF
C25 b0 gnd 0.21fF
C26 vdd a_483_781# 0.22fF
C27 a1 w_238_1377# 0.06fF
C28 w_367_1377# a_350_1365# 0.19fF
C29 a_483_781# a_542_689# 0.02fF
C30 c0 a_396_696# 0.45fF
C31 vdd w_670_905# 0.19fF
C32 a_495_1121# a_518_778# 0.05fF
C33 a3 w_777_1327# 0.06fF
C34 w_559_701# a_483_781# 0.06fF
C35 vdd w_389_701# 0.05fF
C36 a_256_696# w_480_982# 0.06fF
C37 w_670_905# a_685_911# 0.14fF
C38 vdd w_667_821# 0.15fF
C39 a_396_696# w_670_1052# 0.06fF
C40 a_346_1121# a_63_1351# 0.21fF
C41 a_63_1351# a_396_696# 0.58fF
C42 a_396_696# a_685_1058# 0.17fF
C43 a0 a_63_1351# 0.12fF
C44 a_696_771# a_256_696# 0.09fF
C45 a_685_988# a_63_1351# 0.11fF
C46 a_790_1315# w_777_1327# 0.03fF
C47 a_262_689# w_279_701# 0.19fF
C48 a_346_1058# a_116_696# 0.17fF
C49 b0 a_33_1383# 0.21fF
C50 vdd a_130_1315# 0.11fF
C51 b2 a_473_1383# 0.21fF
C52 a_236_1121# w_221_1115# 0.09fF
C53 a_236_1121# gnd 0.08fF
C54 a_256_696# w_331_1115# 0.06fF
C55 c0 a_283_1351# 0.66fF
C56 w_279_701# a_256_696# 0.06fF
C57 w_331_1115# a_369_785# 0.03fF
C58 a_262_689# gnd 0.08fF
C59 vdd w_147_1377# 0.11fF
C60 a_334_788# a_402_689# 0.02fF
C61 a_350_1315# vdd 0.11fF
C62 a_536_696# a_256_696# 0.41fF
C63 a_334_788# a_536_696# 0.09fF
C64 w_331_1052# a_116_696# 0.06fF
C65 b0 w_117_1377# 0.06fF
C66 a_130_1365# a0 0.02fF
C67 w_480_1052# a_256_696# 0.06fF
C68 w_337_1377# b1 0.06fF
C69 a_253_1383# vdd 0.05fF
C70 vdd b0 0.48fF
C71 w_477_821# a_503_1351# 0.06fF
C72 vdd w_337_1327# 0.05fF
C73 a_256_696# gnd 0.85fF
C74 a_283_1351# w_670_1052# 0.06fF
C75 a_334_788# gnd 0.89fF
C76 gnd a_369_785# 0.25fF
C77 w_670_982# vdd 0.18fF
C78 b1 gnd 0.21fF
C79 a_283_1351# a_63_1351# 0.26fF
C80 a_283_1351# a_685_1058# 0.11fF
C81 a_542_778# a_518_778# 0.08fF
C82 a_350_1365# w_337_1377# 0.03fF
C83 a_116_696# a_503_1351# 0.17fF
C84 vdd w_117_1327# 0.05fF
C85 a_262_689# w_249_701# 0.03fF
C86 b2 a2 0.97fF
C87 a_350_1365# gnd 0.08fF
C88 a_122_689# w_109_701# 0.03fF
C89 vdd w_109_701# 0.05fF
C90 a_256_696# w_249_701# 0.06fF
C91 a_790_1365# a3 0.02fF
C92 a_334_788# a_339_785# 0.05fF
C93 a_339_785# a_369_785# 0.08fF
C94 a_732_771# a_696_771# 0.08fF
C95 a_130_1315# w_147_1377# 0.06fF
C96 vdd w_109_651# 0.05fF
C97 a_236_1121# vdd 0.05fF
C98 a_402_639# s2 0.08fF
C99 c0 w_480_982# 0.06fF
C100 w_480_1115# a_396_696# 0.06fF
C101 a_262_689# vdd 0.74fF
C102 w_670_1115# a_685_1121# 0.09fF
C103 a3 a_693_1383# 0.03fF
C104 a_790_1365# a_790_1315# 0.02fF
C105 a_339_785# w_328_821# 0.10fF
C106 gnd a_518_778# 0.34fF
C107 c0 w_139_701# 0.06fF
C108 a_696_771# c0 0.09fF
C109 b0 w_147_1377# 0.06fF
C110 vdd a_256_696# 1.23fF
C111 w_117_1327# a_130_1315# 0.03fF
C112 a_229_792# w_218_821# 0.10fF
C113 a_334_788# vdd 0.22fF
C114 vdd a_369_785# 0.45fF
C115 a_350_1315# w_337_1327# 0.03fF
C116 vdd b1 0.48fF
C117 b2 w_458_1377# 0.06fF
C118 a_732_771# gnd 0.25fF
C119 a_396_696# a_503_1351# 7.17fF
C120 a_536_696# w_670_1115# 0.06fF
C121 a_256_696# a_685_911# 0.08fF
C122 a2 a_570_1315# 0.36fF
C123 a_696_771# a3 0.12fF
C124 a_696_771# a_63_1351# 0.09fF
C125 a_402_689# a_402_639# 0.02fF
C126 a_536_696# c0 0.29fF
C127 vdd a_350_1365# 0.74fF
C128 a_346_1058# a_381_785# 0.05fF
C129 a_256_696# w_670_905# 0.06fF
C130 w_480_1115# a_283_1351# 0.06fF
C131 vdd w_328_821# 0.12fF
C132 c0 w_221_1115# 0.06fF
C133 w_480_1115# a_495_1121# 0.09fF
C134 a3 b3 0.97fF
C135 a_685_1121# a_708_771# 0.05fF
C136 c0 gnd 1.30fF
C137 a_696_771# a_708_771# 1.90fF
C138 a_518_778# a_530_778# 1.15fF
C139 a_63_1351# w_331_1115# 0.06fF
C140 a_402_639# gnd 0.31fF
C141 w_238_1377# a_283_1351# 0.03fF
C142 w_331_1052# a_381_785# 0.03fF
C143 a_536_696# w_670_1052# 0.06fF
C144 a_473_1383# gnd 0.04fF
C145 a_536_696# a_685_1058# 0.03fF
C146 a_536_696# a_63_1351# 0.33fF
C147 a_495_988# a_116_696# 0.08fF
C148 a_495_1058# a_396_696# 0.03fF
C149 w_480_1052# a_63_1351# 0.06fF
C150 a_396_696# w_587_1377# 0.02fF
C151 a_283_1351# a_503_1351# 0.17fF
C152 a_488_778# gnd 0.11fF
C153 gnd a3 0.76fF
C154 gnd a_63_1351# 0.47fF
C155 gnd a_685_1058# 0.08fF
C156 vdd a_518_778# 0.45fF
C157 a_696_771# a_720_771# 0.08fF
C158 a_536_696# a_790_1315# 0.08fF
C159 a_122_639# s0 0.08fF
C160 gnd a_708_771# 0.42fF
C161 a_350_1315# a_256_696# 0.08fF
C162 a_732_771# vdd 0.11fF
C163 b2 w_587_1377# 0.06fF
C164 gnd a_790_1315# 0.31fF
C165 a_122_639# w_139_701# 0.06fF
C166 a2 gnd 0.76fF
C167 a_130_1365# gnd 0.08fF
C168 a2 w_557_1327# 0.06fF
C169 a_229_792# a_224_795# 0.05fF
C170 a_253_1383# b1 0.21fF
C171 w_670_982# a_256_696# 0.06fF
C172 a_350_1315# a_350_1365# 0.02fF
C173 vdd w_670_1115# 0.14fF
C174 a_696_771# a_678_771# 0.70fF
C175 a_696_771# a_744_771# 0.08fF
C176 c4 gnd 0.25fF
C177 a_33_1383# a_63_1351# 0.05fF
C178 a_488_778# a_530_778# 0.08fF
C179 a_122_689# c0 0.02fF
C180 gnd a_720_771# 0.34fF
C181 vdd c0 6.36fF
C182 a2 a_570_1365# 0.02fF
C183 vdd a_402_639# 0.11fF
C184 a1 a_283_1351# 0.12fF
C185 w_218_821# a_259_792# 0.06fF
C186 vdd a_473_1383# 0.05fF
C187 c0 a_685_911# 0.11fF
C188 a_495_988# a_396_696# 0.03fF
C189 a_732_771# w_667_821# 0.06fF
C190 vdd w_670_1052# 0.14fF
C191 vdd a_488_778# 0.11fF
C192 a_122_639# gnd 0.31fF
C193 a_116_696# a_396_696# 0.41fF
C194 vdd a3 0.22fF
C195 a_542_778# a_503_1351# 0.08fF
C196 vdd a_63_1351# 1.05fF
C197 w_807_1377# a3 0.06fF
C198 vdd a_685_1058# 0.16fF
C199 w_18_1377# a0 0.06fF
C200 c0 w_670_905# 0.06fF
C201 a_346_1058# gnd 0.08fF
C202 a_678_771# gnd 0.27fF
C203 gnd a_744_771# 0.17fF
C204 a_685_1121# a_503_1351# 0.21fF
C205 a_696_771# a_503_1351# 0.09fF
C206 vdd a_708_771# 0.11fF
C207 a_488_778# a_483_781# 0.05fF
C208 a_262_689# a_256_696# 0.06fF
C209 w_367_1377# a1 0.06fF
C210 a_130_1365# w_117_1377# 0.03fF
C211 vdd a_790_1315# 0.11fF
C212 a_570_1315# w_587_1377# 0.06fF
C213 w_807_1377# a_790_1315# 0.06fF
C214 vdd a2 0.22fF
C215 a_130_1365# vdd 0.74fF
C216 a_536_696# w_529_701# 0.06fF
C217 w_678_1377# a_693_1383# 0.09fF
C218 a_536_696# a_503_1351# 0.83fF
C219 a_256_696# b1 0.12fF
C220 w_419_701# a_396_696# 0.06fF
C221 c4 vdd 0.20fF
C222 a_732_771# w_670_982# 0.03fF
C223 a_283_1351# a_116_696# 6.72fF
C224 vdd a_720_771# 0.11fF
C225 gnd a_503_1351# 0.38fF
C226 a_350_1365# a_256_696# 0.08fF
C227 a_542_639# w_529_651# 0.03fF
C228 w_667_821# a_708_771# 0.06fF
C229 a_350_1365# b1 0.06fF
C230 a_334_788# w_328_821# 0.03fF
C231 a_369_785# w_328_821# 0.06fF
C232 a_122_689# a_122_639# 0.02fF
C233 a_696_771# w_678_1377# 0.03fF
C234 a_122_639# vdd 0.11fF
C235 a_685_988# a_396_696# 0.17fF
C236 a_229_792# gnd 0.05fF
C237 a_346_1058# vdd 0.16fF
C238 vdd a_678_771# 0.11fF
C239 w_678_1377# b3 0.06fF
C240 vdd a_744_771# 0.13fF
C241 vdd w_389_651# 0.05fF
C242 w_218_821# a_224_795# 0.03fF
C243 a_495_1058# w_480_1052# 0.12fF
C244 c4 w_667_821# 0.03fF
C245 w_667_821# a_720_771# 0.06fF
C246 a_495_1058# gnd 0.08fF
C247 vdd w_458_1377# 0.14fF
C248 a_130_1365# a_130_1315# 0.02fF
C249 a_685_911# a_744_771# 0.05fF
C250 vdd w_480_1115# 0.14fF
C251 b2 a_396_696# 0.12fF
C252 w_670_982# a_63_1351# 0.06fF
C253 vdd w_331_1052# 0.14fF
C254 a_503_1351# a_530_778# 0.08fF
C255 a_130_1365# w_147_1377# 0.19fF
C256 a_495_988# w_480_982# 0.11fF
C257 a_542_778# w_477_821# 0.06fF
C258 vdd w_238_1377# 0.14fF
C259 a1 gnd 0.76fF
C260 w_670_905# a_744_771# 0.03fF
C261 a_495_988# a_542_778# 0.05fF
C262 c0 w_109_651# 0.06fF
C263 a_283_1351# a_396_696# 2.05fF
C264 a_116_696# s0 0.12fF
C265 a_116_696# w_480_982# 0.06fF
C266 a_495_1121# a_396_696# 0.03fF
C267 a_570_1365# w_587_1377# 0.19fF
C268 a_236_1121# c0 0.21fF
C269 a_130_1365# b0 0.06fF
C270 a_542_639# s3 0.08fF
C271 vdd w_529_701# 0.05fF
C272 a_396_696# a_224_795# 0.09fF
C273 vdd a_503_1351# 0.62fF
C274 a_678_771# w_667_821# 0.10fF
C275 w_529_701# a_542_689# 0.03fF
C276 a_116_696# w_139_701# 0.06fF
C277 w_667_821# a_744_771# 0.06fF
C278 a_696_771# a_116_696# 0.09fF
C279 a_495_1058# a_530_778# 0.05fF
C280 c0 a_256_696# 0.61fF
C281 a_334_788# a_402_639# 0.36fF
C282 w_419_701# s2 0.02fF
C283 a_229_792# vdd 0.11fF
C284 a_536_696# a_116_696# 0.25fF
C285 a_495_988# gnd 0.08fF
C286 a_495_1121# a_283_1351# 0.21fF
C287 a_495_1058# vdd 0.16fF
C288 a_256_696# a_63_1351# 3.72fF
C289 w_221_1115# a_116_696# 0.06fF
C290 a_570_1315# a_396_696# 0.08fF
C291 a_283_1351# a_381_785# 0.08fF
C292 vdd w_587_1377# 0.11fF
C293 gnd a_116_696# 0.85fF
C294 a_262_639# s1 0.08fF
C295 s2 a_396_696# 0.12fF
C296 a1 vdd 0.22fF
C297 vdd w_678_1377# 0.14fF
C298 a_396_696# w_480_982# 0.06fF
C299 w_221_1115# a_259_792# 0.03fF
C300 gnd a_259_792# 0.17fF
C301 w_419_701# a_402_689# 0.19fF
C302 a_253_1383# w_238_1377# 0.09fF
C303 a_696_771# a_396_696# 6.93fF
C304 w_477_821# a_530_778# 0.06fF
C305 a_122_639# w_109_651# 0.03fF
C306 a_262_639# a_224_795# 0.36fF
C307 a_346_1121# w_331_1115# 0.09fF
C308 w_18_1377# a_33_1383# 0.09fF
C309 a_224_795# w_249_651# 0.06fF
C310 a_542_639# gnd 0.31fF
C311 a_402_689# a_396_696# 0.06fF
C312 a_488_778# a_518_778# 0.08fF
C313 a_536_696# a_396_696# 3.37fF
C314 vdd w_477_821# 0.14fF
C315 a_685_988# a_536_696# 0.03fF
C316 w_480_1052# a_396_696# 0.06fF
C317 a_495_988# vdd 0.10fF
C318 a_346_1121# gnd 0.08fF
C319 gnd a_396_696# 0.76fF
C320 a_122_689# a_116_696# 0.06fF
C321 a0 gnd 0.76fF
C322 vdd a_116_696# 1.21fF
C323 a_346_1058# a_256_696# 0.03fF
C324 s1 w_279_701# 0.02fF
C325 a_685_988# gnd 0.08fF
C326 w_18_1377# vdd 0.14fF
C327 a_790_1365# w_777_1377# 0.03fF
C328 a_696_771# a_283_1351# 0.09fF
C329 w_477_821# a_483_781# 0.03fF
C330 a_262_639# w_249_651# 0.03fF
C331 a_334_788# w_389_651# 0.06fF
C332 a_116_696# a_685_911# 0.08fF
C333 a1 a_350_1315# 0.36fF
C334 a_732_771# a_708_771# 0.08fF
C335 a_570_1365# a_396_696# 0.08fF
C336 s1 gnd 0.13fF
C337 vdd a_259_792# 0.48fF
C338 w_331_1052# a_256_696# 0.06fF
C339 b2 gnd 0.21fF
C340 a_253_1383# a1 0.03fF
C341 a_116_696# w_670_905# 0.06fF
C342 a1 w_337_1327# 0.06fF
C343 c0 a_63_1351# 6.77fF
C344 a_536_696# a_283_1351# 0.33fF
C345 w_670_1115# a_708_771# 0.03fF
C346 vdd w_218_821# 0.11fF
C347 w_279_701# a_224_795# 0.06fF
C348 w_238_1377# b1 0.06fF
C349 a_536_696# a_224_795# 0.09fF
C350 a_33_1383# a0 0.03fF
C351 vdd w_419_701# 0.11fF
C352 a_283_1351# gnd 0.38fF
C353 b2 a_570_1365# 0.06fF
C354 a_256_696# a_503_1351# 6.82fF
C355 a_732_771# a_720_771# 1.00fF
C356 a_495_1121# gnd 0.08fF
C357 a_790_1365# b3 0.06fF
C358 vdd a_542_639# 0.11fF
C359 w_670_1052# a_685_1058# 0.12fF
C360 gnd a_224_795# 0.80fF
C361 vdd w_777_1327# 0.05fF
C362 gnd a_381_785# 0.17fF
C363 a_542_639# a_542_689# 0.02fF
C364 a_536_696# s3 0.12fF
C365 a_536_696# a_790_1365# 0.08fF
C366 a_696_771# a_693_1383# 0.05fF
C367 a_130_1315# a_116_696# 0.08fF
C368 a_542_639# w_559_701# 0.06fF
C369 a_542_778# w_480_982# 0.03fF
C370 a_262_639# w_279_701# 0.06fF
C371 a_346_1121# vdd 0.05fF
C372 a2 a_473_1383# 0.03fF
C373 vdd a_396_696# 1.09fF
C374 vdd a0 0.22fF
C375 a_542_639# a_483_781# 0.36fF
C376 w_139_701# s0 0.02fF
C377 s3 gnd 0.13fF
C378 gnd a_790_1365# 0.08fF
C379 a_685_988# vdd 0.10fF
C380 a3 a_790_1315# 0.36fF
C381 b3 w_777_1377# 0.06fF
C382 b3 a_693_1383# 0.21fF
C383 a_116_696# w_147_1377# 0.02fF
C384 a_339_785# a_283_1351# 0.37fF
C385 w_480_1115# a_518_778# 0.03fF
C386 vdd w_529_651# 0.05fF
C387 a_396_696# a_685_911# 0.17fF
C388 a_732_771# a_678_771# 0.08fF
C389 a_732_771# a_744_771# 0.52fF
C390 a_262_639# gnd 0.31fF
C391 a_495_1058# a_256_696# 0.17fF
C392 b0 a_116_696# 0.12fF
C393 a_402_689# s2 0.08fF
C394 vdd s1 0.03fF
C395 w_18_1377# b0 0.06fF
C396 w_670_1052# a_720_771# 0.03fF
C397 a_396_696# w_670_905# 0.06fF
C398 b2 vdd 0.48fF
C399 a_122_639# c0 0.36fF
C400 a_570_1315# gnd 0.31fF
C401 a_483_781# w_529_651# 0.06fF
C402 a_570_1315# w_557_1327# 0.03fF
C403 a_685_1058# a_720_771# 0.05fF
C404 gnd a_693_1383# 0.04fF
C405 b2 w_557_1377# 0.06fF
C406 a_396_696# w_389_701# 0.06fF
C407 a_518_778# a_503_1351# 1.59fF
C408 a1 b1 0.97fF
C409 a_346_1058# c0 0.11fF
C410 s2 gnd 0.13fF
C411 a_708_771# a_720_771# 1.45fF
C412 gnd s0 0.13fF
C413 vdd a_283_1351# 0.79fF
C414 a_536_696# a_685_1121# 0.03fF
C415 a_570_1365# a_570_1315# 0.02fF
C416 a_402_639# w_389_651# 0.03fF
C417 a_536_696# a_696_771# 7.08fF
C418 vdd a_495_1121# 0.05fF
C419 a_542_778# gnd 0.17fF
C420 w_109_701# a_116_696# 0.06fF
C421 a1 a_350_1365# 0.02fF
C422 vdd a_224_795# 0.22fF
C423 vdd a_381_785# 0.39fF
C424 w_331_1052# c0 0.06fF
C425 w_458_1377# a_473_1383# 0.09fF
C426 a_685_1121# gnd 0.08fF
C427 a_696_771# gnd 0.47fF
C428 a_536_696# b3 0.12fF
C429 a0 a_130_1315# 0.36fF
C430 w_670_1115# a_503_1351# 0.06fF
C431 vdd s3 0.03fF
C432 a_236_1121# a_116_696# 0.03fF
C433 gnd b3 0.21fF
C434 vdd a_790_1365# 0.74fF
C435 a0 w_147_1377# 0.06fF
C436 a_678_771# a_708_771# 0.08fF
C437 s3 a_542_689# 0.08fF
C438 a_708_771# a_744_771# 0.08fF
C439 w_807_1377# a_790_1365# 0.19fF
C440 c0 a_503_1351# 0.75fF
C441 a_402_689# gnd 0.08fF
C442 a_495_988# a_256_696# 0.17fF
C443 w_367_1377# vdd 0.11fF
C444 a_536_696# gnd 2.96fF
C445 w_559_701# s3 0.02fF
C446 vdd a_262_639# 0.11fF
C447 a_473_1383# a_503_1351# 0.05fF
C448 b0 a0 0.97fF
C449 a_236_1121# a_259_792# 0.05fF
C450 a_256_696# a_116_696# 2.73fF
C451 w_670_982# a_396_696# 0.06fF
C452 vdd w_249_651# 0.05fF
C453 a_542_778# a_530_778# 0.69fF
C454 vdd a_570_1315# 0.11fF
C455 a_685_988# w_670_982# 0.11fF
C456 vdd a_693_1383# 0.05fF
C457 a_488_778# a_503_1351# 0.54fF
C458 vdd w_777_1377# 0.05fF
C459 a0 w_117_1327# 0.06fF
C460 a2 w_458_1377# 0.06fF
C461 c4 a_678_771# 0.05fF
C462 a_63_1351# a_503_1351# 0.17fF
C463 a_678_771# a_720_771# 0.08fF
C464 a_720_771# a_744_771# 0.08fF
C465 vdd s2 0.03fF
C466 a_122_689# s0 0.08fF
C467 vdd s0 0.03fF
C468 vdd w_480_982# 0.18fF
C469 a_570_1365# gnd 0.08fF
C470 a_542_778# vdd 0.30fF
C471 a_122_689# w_139_701# 0.19fF
C472 vdd w_139_701# 0.11fF
C473 vdd a_685_1121# 0.05fF
C474 vdd a_696_771# 0.20fF
C475 a_339_785# gnd 0.10fF
C476 a_253_1383# a_283_1351# 0.05fF
C477 a_229_792# a_63_1351# 0.21fF
C478 a2 a_503_1351# 0.12fF
C479 a_334_788# w_419_701# 0.06fF
C480 w_477_821# a_518_778# 0.06fF
C481 w_480_1052# a_530_778# 0.03fF
C482 a_33_1383# gnd 0.04fF
C483 gnd a_530_778# 0.25fF
C484 a_495_1058# a_63_1351# 0.11fF
C485 vdd b3 0.48fF
C486 vdd w_331_1115# 0.14fF
C487 w_807_1377# b3 0.06fF
C488 vdd a_402_689# 0.74fF
C489 vdd w_279_701# 0.11fF
C490 vdd a_536_696# 0.85fF
C491 w_678_1377# a3 0.06fF
C492 a_346_1121# a_256_696# 0.03fF
C493 a_346_1058# w_331_1052# 0.12fF
C494 w_367_1377# a_350_1315# 0.06fF
C495 w_807_1377# a_536_696# 0.02fF
C496 vdd w_337_1377# 0.05fF
C497 a_536_696# a_542_689# 0.06fF
C498 a_256_696# a_396_696# 3.67fF
C499 a_346_1121# a_369_785# 0.05fF
C500 a_334_788# a_396_696# 0.32fF
C501 vdd w_480_1052# 0.14fF
C502 vdd w_221_1115# 0.14fF
C503 a_685_988# a_256_696# 0.08fF
C504 a_262_689# s1 0.08fF
C505 a_536_696# a_685_911# 0.03fF
C506 a_122_689# gnd 0.08fF
C507 vdd gnd 14.37fF
C508 a_536_696# w_559_701# 0.06fF
C509 vdd w_557_1327# 0.05fF
C510 gnd a_542_689# 0.08fF
C511 a_696_771# w_667_821# 0.06fF
C512 a_536_696# a_483_781# 0.32fF
C513 a2 w_587_1377# 0.06fF
C514 gnd a_685_911# 0.08fF
C515 a_536_696# w_670_905# 0.06fF
C516 s1 a_256_696# 0.12fF
C517 a_402_689# w_389_701# 0.03fF
C518 a_495_988# c0 0.11fF
C519 vdd a_570_1365# 0.74fF
C520 a_483_781# gnd 0.89fF
C521 a_570_1365# w_557_1377# 0.03fF
C522 w_458_1377# a_503_1351# 0.03fF
C523 c0 a_116_696# 6.02fF
C524 a_262_689# a_224_795# 0.02fF
C525 vdd w_249_701# 0.05fF
C526 a_339_785# vdd 0.11fF
C527 w_477_821# a_488_778# 0.10fF
C528 a_256_696# a_283_1351# 7.28fF
C529 a_283_1351# a_369_785# 1.29fF
C530 vdd a_33_1383# 0.05fF
C531 a_256_696# a_224_795# 0.33fF
C532 vdd a_530_778# 0.37fF
C533 s3 Gnd 1.08fF
C534 a_542_639# Gnd 1.09fF
C535 a_542_689# Gnd 0.88fF
C536 s2 Gnd 1.08fF
C537 a_402_639# Gnd 1.09fF
C538 a_402_689# Gnd 0.88fF
C539 s1 Gnd 1.08fF
C540 a_262_639# Gnd 1.09fF
C541 a_262_689# Gnd 0.88fF
C542 s0 Gnd 1.08fF
C543 a_122_639# Gnd 1.09fF
C544 a_122_689# Gnd 0.88fF
C545 c4 Gnd 2.29fF
C546 a_483_781# Gnd 3.25fF
C547 a_334_788# Gnd 3.30fF
C548 a_224_795# Gnd 3.01fF
C549 a_678_771# Gnd 0.63fF
C550 a_488_778# Gnd 0.52fF
C551 a_339_785# Gnd 0.43fF
C552 a_229_792# Gnd 0.32fF
C553 a_744_771# Gnd 1.30fF
C554 a_685_911# Gnd 0.61fF
C555 a_732_771# Gnd 2.34fF
C556 a_542_778# Gnd 2.05fF
C557 a_685_988# Gnd 0.51fF
C558 a_495_988# Gnd 0.51fF
C559 a_720_771# Gnd 3.29fF
C560 a_530_778# Gnd 2.95fF
C561 a_381_785# Gnd 2.74fF
C562 a_685_1058# Gnd 0.42fF
C563 a_495_1058# Gnd 0.42fF
C564 a_346_1058# Gnd 0.42fF
C565 a_708_771# Gnd 4.17fF
C566 a_518_778# Gnd 3.79fF
C567 a_369_785# Gnd 3.58fF
C568 a_259_792# Gnd 3.38fF
C569 a_685_1121# Gnd 0.32fF
C570 a_495_1121# Gnd 0.32fF
C571 a_346_1121# Gnd 0.32fF
C572 a_236_1121# Gnd 0.32fF
C573 c0 Gnd 18.74fF
C574 a_536_696# Gnd 21.08fF
C575 a_696_771# Gnd 15.60fF
C576 a_790_1315# Gnd 1.09fF
C577 a_693_1383# Gnd 0.32fF
C578 b3 Gnd 3.91fF
C579 a3 Gnd 3.51fF
C580 a_790_1365# Gnd 0.88fF
C581 a_396_696# Gnd 21.46fF
C582 a_503_1351# Gnd 14.24fF
C583 a_570_1315# Gnd 1.09fF
C584 a_473_1383# Gnd 0.32fF
C585 b2 Gnd 3.91fF
C586 a2 Gnd 3.51fF
C587 a_570_1365# Gnd 0.88fF
C588 a_256_696# Gnd 20.55fF
C589 a_283_1351# Gnd 13.67fF
C590 a_350_1315# Gnd 1.09fF
C591 a_253_1383# Gnd 0.32fF
C592 b1 Gnd 3.91fF
C593 a1 Gnd 3.51fF
C594 a_350_1365# Gnd 0.88fF
C595 gnd Gnd 27.15fF
C596 a_116_696# Gnd 18.02fF
C597 a_63_1351# Gnd 13.77fF
C598 vdd Gnd 24.27fF
C599 a_130_1315# Gnd 1.09fF
C600 a_33_1383# Gnd 0.32fF
C601 b0 Gnd 3.91fF
C602 a0 Gnd 3.51fF
C603 a_130_1365# Gnd 0.88fF
C604 w_529_651# Gnd 0.48fF
C605 w_389_651# Gnd 0.48fF
C606 w_249_651# Gnd 0.48fF
C607 w_109_651# Gnd 0.48fF
C608 w_559_701# Gnd 1.12fF
C609 w_529_701# Gnd 0.48fF
C610 w_419_701# Gnd 1.12fF
C611 w_389_701# Gnd 0.48fF
C612 w_279_701# Gnd 1.12fF
C613 w_249_701# Gnd 0.48fF
C614 w_139_701# Gnd 1.12fF
C615 w_109_701# Gnd 0.48fF
C616 w_667_821# Gnd 1.85fF
C617 w_477_821# Gnd 1.61fF
C618 w_328_821# Gnd 1.37fF
C619 w_218_821# Gnd 1.12fF
C620 w_670_905# Gnd 1.85fF
C621 w_670_982# Gnd 1.61fF
C622 w_480_982# Gnd 1.61fF
C623 w_670_1052# Gnd 1.37fF
C624 w_480_1052# Gnd 1.37fF
C625 w_331_1052# Gnd 1.37fF
C626 w_670_1115# Gnd 1.12fF
C627 w_480_1115# Gnd 1.12fF
C628 w_331_1115# Gnd 1.12fF
C629 w_221_1115# Gnd 1.12fF
C630 w_777_1327# Gnd 0.48fF
C631 w_557_1327# Gnd 0.48fF
C632 w_337_1327# Gnd 0.48fF
C633 w_117_1327# Gnd 0.48fF
C634 w_807_1377# Gnd 1.12fF
C635 w_777_1377# Gnd 0.48fF
C636 w_678_1377# Gnd 1.12fF
C637 w_587_1377# Gnd 1.12fF
C638 w_557_1377# Gnd 0.48fF
C639 w_458_1377# Gnd 1.12fF
C640 w_367_1377# Gnd 1.12fF
C641 w_337_1377# Gnd 0.48fF
C642 w_238_1377# Gnd 1.12fF
C643 w_147_1377# Gnd 1.12fF
C644 w_117_1377# Gnd 0.48fF
C645 w_18_1377# Gnd 1.12fF


.tran 1n 20n

.control
set hcopypscolor=1
set color0=white
set color1=black
run
set curplottitle="jal_2023102066_adder"

meas tran worst_case_delay trig v(A0) val=0.9 fall=1 targ v(S2) val=0.9 fall=1

plot v(c0)
plot a0 a1+2 a2+4 a3+6
plot b0 b1+2 b2+4 b3+6
plot s0 s1+2 s2+4 s3+6 c4+8
.endc

.end